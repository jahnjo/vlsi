* Component: $VLSI/Project/test  Viewpoint: default
.INCLUDE $VLSI/Project/test/default/test_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 150N

* --- Waveform Outputs
.PROBE TRAN V(ENABLE)
.PROBE TRAN V(CLK)
.PROBE TRAN V(A)
.PROBE TRAN V(B)
.PROBE TRAN V(X)
.PROBE TRAN V(Y)

* --- Params
.TEMP 27

* --- Forces
VFORCE__A A GROUND PULSE (0 2.5v 15n 1n 1n 20n 40n)
VFORCE__B B GROUND PULSE (0 2.5v 35n 1n 1n 40n 80n)
VFORCE__Enable ENABLE GROUND dc 2.5v
VFORCE__Enable_1 CLK GROUND PULSE (0 2.5v 0n 1n 1n 10n 20n)
VFORCE__Enable_2 VDD GROUND dc 2.5v

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

