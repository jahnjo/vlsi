* Component: $VLSI/Project/inv  Viewpoint: default
.INCLUDE $VLSI/Project/inv/default/inv_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 100N

* --- Waveform Outputs
.PROBE TRAN V(IN)
.PROBE TRAN V(VDD)
.PROBE TRAN V(OUT)

* --- Params
.TEMP 27

* --- Forces
VFORCE___VDD VDD GROUND dc 2.5v
VFORCE__IN IN GROUND PULSE (0 2.5v 25n 1n 1n 25n 50n)

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

