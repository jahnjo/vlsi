*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'egrvlsi07' on Thu Apr  4 2019 at 15:46:07

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $VLSI/Project/Mux21
*
.subckt MUX21  Y A B S

        M6 Y N$46 A GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p ps=1.28u
+  pd=1.28u
        M3 Y S A VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M5 Y S B GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p ps=1.28u
+  pd=1.28u
        M4 Y N$46 B VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M2 N$46 S VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M1 N$46 S GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
.ends MUX21

*
* Component pathname : $VLSI/Project/Mux41
*
.subckt MUX41  OUT1 IN0 IN1 IN2 IN3 S0 S1

        X_MUX213 OUT1 N$2 N$4 S1 MUX21
        X_MUX212 N$4 IN2 IN3 S0 MUX21
        X_MUX211 N$2 IN0 IN1 S0 MUX21
.ends MUX41

*
* Component pathname : $VLSI/Project/inv
*
.subckt INV  OUT IN

        M2 OUT IN VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M1 OUT IN GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
.ends INV

*
* Component pathname : $VLSI/Project/or
*
.subckt OR  Y A B

        M6 Y N$22 GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M5 Y N$22 VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M4 N$22 A GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M3 N$22 B GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M2 N$22 B N$13 VDD pmos w=2.7u l=0.13u m=1 as=0.918p ad=0.918p ps=3.38u
+  pd=3.38u
        M1 N$13 A VDD VDD pmos w=2.7u l=0.13u m=1 as=0.918p ad=0.918p ps=3.38u
+  pd=3.38u
.ends OR

*
* Component pathname : $VLSI/Project/and
*
.subckt AND  Y A B

        M6 Y N$54 GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M5 Y N$54 VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M4 N$54 B VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M3 N$54 A VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M2 N$29 B GROUND GROUND nmos w=1.2u l=0.13u m=1 as=0.408p ad=0.408p
+  ps=1.88u pd=1.88u
        M1 N$54 A N$29 GROUND nmos w=1.2u l=0.13u m=1 as=0.408p ad=0.408p
+  ps=1.88u pd=1.88u
.ends AND

*
* Component pathname : $VLSI/Project/Adder
*
.subckt ADDER  COUT S A B CIN

        M18 N$145 CIN N$165 GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M17 N$145 CIN N$159 VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M16 N$159 B N$157 VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M15 N$157 A VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M24 N$47 CIN GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M23 N$47 B GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M22 N$47 A GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M21 N$145 N$210 N$47 GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M14 N$145 N$210 N$37 VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M13 N$37 CIN VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M12 N$37 B VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M11 N$37 A VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M10 N$7 B VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M9 N$10 B VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M8 N$10 A VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M7 N$210 A N$7 VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M6 N$210 A N$19 GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M5 N$210 CIN N$14 GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M4 N$19 B GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M3 N$14 B GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M2 N$210 CIN N$10 VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M1 N$14 A GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M28 S N$145 GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M27 S N$145 VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M26 COUT N$210 GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M25 COUT N$210 VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M20 N$167 A GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
        M19 N$165 B N$167 GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
.ends ADDER

*
* MAIN CELL: Component pathname : $VLSI/Project/alu
*
        X_MUX411 RESULT N$32 N$32 N$31 N$30 ALUOP_0 ALUOP_1 MUX41
        X_INV N$41 B INV
        X_B_MUX N$44 B N$41 ALUOP_0 MUX21
        X_OR N$30 A B OR
        X_AND N$31 A B AND
        X_ADD_SUB COUT N$32 A N$44 ALUOP_0 ADDER
*
.end
