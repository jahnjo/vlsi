*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'egrvlsi07' on Mon Apr  8 2019 at 17:02:25

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $VLSI/Project/and
*
.subckt AND  Y A B

        M6 Y N$54 GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M5 Y N$54 VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M4 N$54 B VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M3 N$54 A VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M2 N$29 B GROUND GROUND nmos w=1.2u l=0.13u m=1 as=0.408p ad=0.408p
+  ps=1.88u pd=1.88u
        M1 N$54 A N$29 GROUND nmos w=1.2u l=0.13u m=1 as=0.408p ad=0.408p
+  ps=1.88u pd=1.88u
.ends AND

*
* Component pathname : $VLSI/Project/and3
*
.subckt AND3  Y A B C

        X_AND2 Y N$10 C AND
        X_AND1 N$10 A B AND
.ends AND3

*
* Component pathname : $VLSI/Project/inv
*
.subckt INV  OUT IN

        M2 OUT IN VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M1 OUT IN GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
.ends INV

*
* MAIN CELL: Component pathname : $VLSI/Project/decoder
*
        X_AND38 REG7 RD_0 RD_1 RD_2 AND3
        X_AND37 REG6 N$31 RD_1 RD_2 AND3
        X_AND36 REG5 RD_0 N$45 RD_2 AND3
        X_AND35 REG4 N$31 N$45 RD_2 AND3
        X_AND34 REG3 RD_0 RD_1 N$51 AND3
        X_AND33 REG2 N$31 RD_1 N$51 AND3
        X_AND32 REG1 RD_0 N$45 N$51 AND3
        X_AND31 REG0 N$31 N$45 N$51 AND3
        X_INV3 RD_0 N$31 INV
        X_INV2 RD_1 N$45 INV
        X_INV1 RD_2 N$51 INV
*
.end
