* Component: $VLSI/Project/DFF  Viewpoint: default
.INCLUDE $VLSI/Project/DFF/default/DFF_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 100N

* --- Waveform Outputs
.PROBE TRAN V(CLK)
.PROBE TRAN V(D)
.PROBE TRAN V(Q)
.PROBE TRAN V(Q_BAR)

* --- Params
.TEMP 27
.PARAM t_sweep=0 
.STEP PARAM t_sweep 0n 100n INCR 1n

* --- Forces
VFORCE__D D GROUND PULSE (0 2.5v 25n 1n 1n 25n 50n)
VFORCE__CLK CLK GROUND PULSE (0 2.5v 10n 1n 1n 10n 20n)
VFORCE___VDD VDD GROUND dc 2.5v

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

