* Component: $VLSI/Project/Mux21  Viewpoint: default
.INCLUDE $VLSI/Project/Mux21/default/Mux21_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 100N

* --- Waveform Outputs
.PROBE TRAN V(S)
.PROBE TRAN V(A)
.PROBE TRAN V(B)
.PROBE TRAN V(Y)

* --- Params
.TEMP 27
.PARAM t_sweep=0 
.STEP PARAM t_sweep 0n 100n INCR 1n

* --- Forces
VFORCE___VDD VDD GROUND dc 2.5v
VFORCE__A A GROUND PULSE (0 2.5 0n 1n 1n 100n 100n)
VFORCE__B B GROUND PULSE (0 2.5 0n 1n 1n 100n 100n)
VFORCE__S S GROUND PULSE (0 2.5 25n 1n 1n 25n 50n)

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

