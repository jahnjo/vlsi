* Component: $VLSI/Project/DFFen  Viewpoint: default
.INCLUDE $VLSI/Project/DFFen/default/DFFen_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 500N

* --- Waveform Outputs
.PROBE TRAN V(D)
.PROBE TRAN V(EN)
.PROBE TRAN V(CLK)
.PROBE TRAN V(Q)

* --- Params
.TEMP 27

* --- Forces
VFORCE__D D GROUND PULSE (0 2.5v 20n 1n 1n 30n 60n)
VFORCE__En EN GROUND PULSE (0 2.5v 25n 1n 1n 100n 200n)
VFORCE__CLK CLK GROUND PULSE (0 2.5v 15n 1n 1n 15n 30n)
VFORCE___VDD VDD GROUND dc 2.5v

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

