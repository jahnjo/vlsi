* Component: $VLSI/Project/reg  Viewpoint: default
.INCLUDE $VLSI/Project/reg/default/reg_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 400N

* --- Waveform Outputs
.PROBE TRAN V(BUSW)
.PROBE TRAN V(CLK)
.PROBE TRAN V(REG_W)
.PROBE TRAN V(DEC0)
.PROBE TRAN V(DEC1)
.PROBE TRAN V(DEC2)
.PROBE TRAN V(DEC3)
.PROBE TRAN V(DEC4)
.PROBE TRAN V(DEC5)
.PROBE TRAN V(DEC6)
.PROBE TRAN V(DEC7)
.PROBE TRAN V(RT0)
.PROBE TRAN V(RT1)
.PROBE TRAN V(RT2)
.PROBE TRAN V(RS0)
.PROBE TRAN V(RS1)
.PROBE TRAN V(RS2)
.PROBE TRAN V(BUSA)
.PROBE TRAN V(BUSB)

* --- Params
.TEMP 27

* --- Forces
VFORCE__BusW BUSW GROUND PULSE (0 2.5v 0 1n 1n 100n 200n)
VFORCE__clk CLK GROUND PULSE (0 2.5v 0 1n 1n 10n 20n)
VFORCE__Reg_W REG_W GROUND PULSE (0 2.5v 0 1n 1n 400n 800n)
VFORCE__dec0 DEC0 GROUND PULSE (0 2.5v 0 1n 1n 20n 400n)
VFORCE__dec1 DEC1 GROUND PULSE (0 2.5v 20n 1n 1n 20n 400n)
VFORCE__dec2 DEC2 GROUND PULSE (0 2.5v 40n 1n 1n 20n 400n)
VFORCE__dec3 DEC3 GROUND PULSE (0 2.5v 60n 1n 1n 20n 400n)
VFORCE__dec4 DEC4 GROUND PULSE (0 2.5v 80n 1n 1n 20n 400n)
VFORCE__dec5 DEC5 GROUND PULSE (0 2.5v 100n 1n 1n 20n 400n)
VFORCE__dec6 DEC6 GROUND PULSE (0 2.5v 120n 1n 1n 20n 400n)
VFORCE__dec7 DEC7 GROUND PULSE (0 2.5v 140n 1n 1n 20n 400n)
VFORCE__Rt0 RT0 GROUND PULSE (0 2.5v 40n 1n 1n 20n 40n)
VFORCE__Rt1 RT1 GROUND PULSE (0 2.5v 60n 1n 1n 40n 80n)
VFORCE__Rt2 RT2 GROUND PULSE (0 2.5v 100n 1n 1n 80n 160n)
VFORCE__Rs0 RS0 GROUND PULSE (0 2.5v 40n 1n 1n 20n 40n)
VFORCE__Rs1 RS1 GROUND PULSE (0 2.5v 60n 1n 1n 40n 80n)
VFORCE__Rs2 RS2 GROUND PULSE (0 2.5v 100n 1n 1n 80n 160n)
VFORCE___VDD VDD GROUND dc 1

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

