*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'egrvlsi07' on Wed Mar 27 2019 at 13:25:02

*
* Globals.
*
.global GROUND VDD

*
* MAIN CELL: Component pathname : $VLSI/Project/Mux21
*
        M6 Y N$46 A GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M3 Y S A VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u pd=2.68u
        M5 Y S B GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M4 Y N$46 B VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M2 N$46 S VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M1 N$46 S GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
*
.end
