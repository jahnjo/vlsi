*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'egrvlsi07' on Tue Mar 26 2019 at 17:04:21

*
* Globals.
*
.global VDD GROUND

*
* MAIN CELL: Component pathname : $VLSI/Project/Mux21
*
        M6 A N$46 Y N$55 nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M3 A S Y N$56 pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u pd=2.68u
        M5 B S Y N$57 nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u pd=2.68u
        M4 B N$46 Y N$62 pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M2 N$46 S VDD VDD pmos w=2u l=0.13u m=1 as=0.68p ad=0.68p ps=2.68u
+  pd=2.68u
        M1 N$46 S GROUND GROUND nmos w=2u l=0.13u m=1 as=0.68p ad=0.68p
+  ps=2.68u pd=2.68u
*
.end
