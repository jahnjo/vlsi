* Component: $VLSI/Project/imm_mux  Viewpoint: default
.INCLUDE $VLSI/Project/imm_mux/default/imm_mux_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 100N

* --- Waveform Outputs
.PROBE TRAN V(INPUT_SELECT)
.PROBE TRAN V(RESULT_3)
.PROBE TRAN V(RESULT_2)
.PROBE TRAN V(RESULT_1)
.PROBE TRAN V(RESULT_0)
.PROBE TRAN V(IMM_3)
.PROBE TRAN V(IMM_2)
.PROBE TRAN V(IMM_1)
.PROBE TRAN V(IMM_0)
.PROBE TRAN V(BUSW_RESULT_3)
.PROBE TRAN V(BUSW_RESULT_2)
.PROBE TRAN V(BUSW_RESULT_1)
.PROBE TRAN V(BUSW_RESULT_0)

* --- Params
.TEMP 27

* --- Forces
VFORCE__input_select INPUT_SELECT GROUND PULSE (0 2.5v 0 1n 1n 50n 100n)
VFORCE__result RESULT_3 GROUND PULSE (0 2.5v 100n 1n 1n 50n 100n)
VFORCE__result_1 RESULT_2 GROUND PULSE (0 2.5v 100n 1n 1n 50n 100n)
VFORCE__result_2 RESULT_1 GROUND PULSE (0 2.5v 100n 1n 1n 50n 100n)
VFORCE__result_3 RESULT_0 GROUND PULSE (0 2.5v 100n 1n 1n 50n 100n)
VFORCE__imm IMM_3 GROUND PULSE (0 2.5v 0n 1n 1n 100n 200n)
VFORCE__imm_1 IMM_2 GROUND PULSE (0 2.5v 0n 1n 1n 100n 200n)
VFORCE__imm_2 IMM_1 GROUND PULSE (0 2.5v 0n 1n 1n 100n 200n)
VFORCE__imm_3 IMM_0 GROUND PULSE (0 2.5v 0n 1n 1n 100n 200n)
VFORCE___VDD VDD GROUND dc 2.5v

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

