*
* .CONNECT statements
*
.CONNECT GROUND 0


* ELDO netlist generated with ICnet by 'egrvlsi07' on Wed Apr 17 2019 at 13:25:07

*
* Globals.
*
.global VDD GROUND

*
* Component pathname : $VLSI/Project/or
*
.subckt OR  Y A B

        M6 Y N$22 GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M5 Y N$22 VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M4 N$22 A GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M3 N$22 B GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M2 N$22 B N$13 VDD pmos w=2.7u l=0.13u m=1 as=0.918p ad=0.918p ps=3.38u
+  pd=3.38u
        M1 N$13 A VDD VDD pmos w=2.7u l=0.13u m=1 as=0.918p ad=0.918p ps=3.38u
+  pd=3.38u
.ends OR

*
* Component pathname : $VLSI/Project/or3
*
.subckt OR3  Y A B C

        X_OR2 Y N$5 C OR
        X_OR1 N$5 A B OR
.ends OR3

*
* Component pathname : $VLSI/Project/and
*
.subckt AND  Y A B

        M6 Y N$54 GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
        M5 Y N$54 VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M4 N$54 B VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M3 N$54 A VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M2 N$29 B GROUND GROUND nmos w=1.2u l=0.13u m=1 as=0.408p ad=0.408p
+  ps=1.88u pd=1.88u
        M1 N$54 A N$29 GROUND nmos w=1.2u l=0.13u m=1 as=0.408p ad=0.408p
+  ps=1.88u pd=1.88u
.ends AND

*
* Component pathname : $VLSI/Project/and3
*
.subckt AND3  Y A B C

        X_AND2 Y N$10 C AND
        X_AND1 N$10 A B AND
.ends AND3

*
* Component pathname : $VLSI/Project/inv
*
.subckt INV  OUT IN

        M2 OUT IN VDD VDD pmos w=1.35u l=0.13u m=1 as=0.459p ad=0.459p ps=2.03u
+  pd=2.03u
        M1 OUT IN GROUND GROUND nmos w=0.6u l=0.13u m=1 as=0.204p ad=0.204p
+  ps=1.28u pd=1.28u
.ends INV

*
* MAIN CELL: Component pathname : $VLSI/Project/control
*
        X_OR35 ALU_SRC N$41 N$48 PC_SRC OR3
        X_OR3 ALU_OP_0 N$59 PC_SRC OR
        X_OR34 N$59 N$35 N$56 N$48 OR3
        X_OR2 ALU_OP_1 N$53 N$48 OR
        X_OR33 N$53 N$37 N$41 N$56 OR3
        X_OR1 REG_WRITE N$46 N$48 OR
        X_OR32 N$46 N$39 N$41 N$56 OR3
        X_OR31 N$39 N$33 N$35 N$37 OR3
        X_BEQ PC_SRC N$30 OP_1 OP_2 AND3
        X_ORI N$48 OP_0 N$27 OP_2 AND3
        X_OR N$56 N$30 N$27 OP_2 AND3
        X_ANDI N$41 OP_0 OP_1 N$20 AND3
        X_AND N$37 N$30 OP_1 N$20 AND3
        X_SUB N$35 OP_0 N$27 N$20 AND3
        X_ADD N$33 N$30 N$27 N$20 AND3
        X_INV3 N$30 OP_0 INV
        X_INV2 N$27 OP_1 INV
        X_INV1 N$20 OP_2 INV
*
.end
