* Component: $VLSI/Project/alu  Viewpoint: default
.INCLUDE $VLSI/Project/alu/default/alu_default.spi
.INCLUDE $GENERIC13/models/include_all
.OPTION NOASCII
.OPTION MODWL
.OPTION ENGNOT
.OPTION AEX

* --- Singles

* - Analysis Setup - Trans
.TRAN 0 500N

* --- Waveform Outputs
.PROBE TRAN V(ALUOP_1)
.PROBE TRAN V(ALUOP_0)
.PROBE TRAN V(A)
.PROBE TRAN V(B)
.PROBE TRAN V(RESULT)
.PROBE TRAN V(COUT)

* --- Params
.TEMP 27

* --- Forces
VFORCE__A A GROUND PULSE (0 2.5v 0 1n 1n 500n 1000n)
VFORCE__B B GROUND PULSE (0 2.5v 0 1n 1n 25n 50n)
VFORCE__ALUop ALUOP_0 GROUND PULSE (0 2.5v 100n 1n 1n 50n 100n)
VFORCE__ALUop_1 ALUOP_1 GROUND PULSE (0 2.5v 200n 1n 1n 200n 400n)
VFORCE__ALUop_2 VDD GROUND dc 2.5v

* --- Libsetup
.LIB key=MOS $GENERIC13/models/lib.eldo TT
.LIB key=MOS_33 $GENERIC13/models/lib.eldo TT_33
.LIB key=MOS_lvt $GENERIC13/models/lib.eldo TT_lvt
.LIB key=MOS_hvt $GENERIC13/models/lib.eldo TT_hvt
.LIB key=BIP $GENERIC13/models/lib.eldo TT_BIP
.LIB key=BIP_NPN $GENERIC13/models/lib.eldo TT_BIP_NPN
.LIB key=RES $GENERIC13/models/lib.eldo TT_RES

